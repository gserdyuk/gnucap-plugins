A 5-R noise circuit
*
*  +- R1-+--R3--+----
*  |     |      |    |
*  V     R2     R4  RL
*  |     |      |    | 
* ---   ---    ---  ---
*

.subckt res4 in out
R1  in 12  100
R2  12 0   50.K
R3  12 out 500
R4  out 0 10.K
.ends

Vin 1 0 ac 1 dc 0

*X1  1 3 res4
R1  1 12  100
R2  12 0   50.K
R3  12 3 500
R4  3 0 10.K

RL  3 0 5.K

.noise v(3) vin dec 1 10. 100 
.end
