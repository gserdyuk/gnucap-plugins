A 5-R noise circuit
*
*  +- C1-+--C2--+----
*  |     |      |    |
*  V     R2     R4  RL
*  |     |      |    | 
* ---   ---    ---  ---
*
.subckt res4 in out
C1  in 2  20u
R2  2 0   50.K
C3  2 out 4u
R4  out 0 10.K
.ends

Vin 1 0 ac 1 dc 0
X1  1 3 res4
RL  3 0 5.K

.print noise all
.noise v(3) vin dec 2 10. 1000
.end
