A 5-R noise circuit
*
*  +- R1-+---
*  |         |
*  V         RL
*  |         | 
* ---       ---
*
.subckt res_sub in out
R1  in out 100
.ends

Vin 1 0 ac 1 dc 0
X1  1 3 res_sub
RL  3 0 5.K

.noise v(3) vin dec 1 10. 100 
.end
